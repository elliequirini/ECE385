module color_table(input [7:0] color,
						 output logic [7:0]  Red, Green, Blue);


						 
endmodule