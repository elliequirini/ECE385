module BouncingBall();

endmodule