module LC3_Processor();