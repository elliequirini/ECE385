module testbench ();

endmodule